module ansi_module_b (
  input logic hej
);

  logic a;
  logic b;

endmodule
